module register_MEM_WB(
    input [3:0] opcode
);

endmodule