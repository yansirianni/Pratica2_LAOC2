module memoryAccess();

endmodule