module instructionExecute_Control(
    
);

endmodule // instructionExecute_Control