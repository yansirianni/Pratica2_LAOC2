module register_IF_ID(
    input [3:0] opcode
);

endmodule