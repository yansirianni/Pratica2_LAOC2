module writeBack();

endmodule