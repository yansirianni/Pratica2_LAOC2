module instructionDecode_Control();

endmodule // instructionDecode_Control