module register_IF_ID(
    input [3:0] opcode;
	 input [19:0] instruction;
	 output [19:0] data_out;
);

endmodule