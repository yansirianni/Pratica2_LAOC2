module register_EX_MEM(
    input [3:0] opcode
);

endmodule