module register_ID_EX(
    input [3:0] opcode
);

endmodule