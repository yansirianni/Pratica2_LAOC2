module instructionFetch();

endmodule