module instructionDecode();

endmodule