module memoryAccess(address, out);
    input [19:0] address;
    output [19:0] out;

    assign out = address; 
endmodule