module register_MEM_WB();

endmodule