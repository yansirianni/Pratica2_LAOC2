module memoryAccess_Control(
    
);

endmodule // memoryAccess_Control