module instructionDecode_Control(clock,reset,opcode_in,);

    always @() begin
        
    end

endmodule // instructionDecode_Control