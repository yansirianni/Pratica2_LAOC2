module instructionFetch();

//Automático

endmodule