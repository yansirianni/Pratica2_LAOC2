module instructionExecute();

endmodule