module register_EX_MEM();

endmodule