module instructionDecode();

endmodule

