module writeBack_Control(
    
);

endmodule // writeBack_Control