module register_IF_ID();

endmodule